`define INWD4
// `define INWD6
// `define INWD8
// `define INWD10


`define INWD 4
`define LOGINWD 2
`define CNTWD `INWD
