// `define INWD4
// `define INWD6
`define INWD8
// `define INWD10


`define INWD 8
`define LOGINWD 3
`define CNTWD `INWD
